magic
tech scmos
timestamp 1594232584
<< nwell >>
rect -24 -9 28 26
<< ntransistor >>
rect -8 -39 -5 -29
rect 6 -39 9 -29
<< ptransistor >>
rect -8 0 -5 18
rect 6 0 9 18
<< ndiffusion >>
rect -11 -34 -8 -29
rect -16 -39 -8 -34
rect -5 -39 6 -29
rect 9 -34 15 -29
rect 9 -39 20 -34
<< pdiffusion >>
rect -11 13 -8 18
rect -16 0 -8 13
rect -5 13 -2 18
rect 3 13 6 18
rect -5 0 6 13
rect 9 13 15 18
rect 9 0 20 13
<< ndcontact >>
rect -16 -34 -11 -29
rect 15 -34 20 -29
<< pdcontact >>
rect -16 13 -11 18
rect -2 13 3 18
rect 15 13 20 18
<< polysilicon >>
rect -8 18 -5 22
rect 6 18 9 22
rect -8 -12 -5 0
rect -8 -29 -5 -17
rect 6 -20 9 0
rect 6 -29 9 -25
rect -8 -41 -5 -39
rect 6 -41 9 -39
<< polycontact >>
rect -10 -17 -5 -12
rect 4 -25 9 -20
<< metal1 >>
rect -16 26 20 30
rect -16 18 -11 26
rect 15 18 20 26
rect -2 -12 3 13
rect -13 -17 -10 -12
rect -2 -16 20 -12
rect -13 -25 4 -20
rect 15 -29 20 -16
<< labels >>
rlabel pdcontact -14 17 -14 17 1 VDD!
rlabel metal1 -13 -17 -13 -12 1 va
rlabel metal1 -13 -25 -13 -20 1 vb
rlabel metal1 20 -16 20 -12 1 vout
rlabel ndcontact -14 -30 -14 -30 1 GND!
<< end >>
